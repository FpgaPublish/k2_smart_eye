// --------------------------------------------------------------------
// interface
`include "./lib_interface/data_interface.sv"
// --------------------------------------------------------------------
// VIP
`include "./lib_vip/vip_read_imag.sv"
// --------------------------------------------------------------------
// phase
`include "./lib_phase/file_phase.sv"
// --------------------------------------------------------------------
// main phase
`include "./lib_phase/main_phase.sv"

