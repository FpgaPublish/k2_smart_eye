// --------------------------------------------------------------------
// imag info
`define NB_IMAG_W 480
`define NB_IMAG_H 320
// --------------------------------------------------------------------
// clock time
`define NB_SYS_PER #10
