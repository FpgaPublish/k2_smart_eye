/****************************************************************
 * File : versal_cips_ps_vip_v1_0_5_unused_ports.sv
 *
 * Date : 2015-16
 *
 * Description : Default value driving for unused ports.
 *
 *****************************************************************************/

//////////////////////Everest Unused Ports////////////////////////////

////////////////////////Versal CIPS PS VIP Unused Ports////////////////////////////
  assign   	ADMA2PLCACK = 0;
  assign   	ADMA2PLTVLD = 0;
  assign 	CCI_NOC_0 = 0;
  assign 	CCI_NOC_1 = 0;
  assign 	CCI_NOC_2 = 0;
  assign 	CCI_NOC_3 = 0;
  assign 	CFUEOS = 0;
//  assign 	CPMOSCCLKDIV2 = 0;  // CR-1097551
  assign 	EMIOCAN0PHYTX = 0;
  assign 	EMIOCAN1PHYTX = 0;
  assign   	EMIOENET0DMABUSWIDTH = 0;
  assign 	EMIOENET0DMATXENDTOG = 0;
  assign   	EMIOENET0GEMTSUTIMERCNT = 0;
  assign   	EMIOENET0GMIITXD = 0;
  assign 	EMIOENET0GMIITXEN = 0;
  assign 	EMIOENET0GMIITXER = 0;
  assign 	EMIOENET0MDIOMDC = 0;
  assign 	EMIOENET0MDIOO = 0;
  assign 	EMIOENET0MDIOTN = 0;
  assign 	EMIOENET0RXWDATA = 0;
  assign 	EMIOENET0RXWEOP = 0;
  assign 	EMIOENET0RXWERR = 0;
  assign 	EMIOENET0RXWFLUSH = 0;
  assign 	EMIOENET0RXWSOP = 0;
  assign 	EMIOENET0RXWSTATUS = 0;
  assign 	EMIOENET0RXWWR = 0;
  assign 	EMIOENET0SPEEDMODE = 0;
  assign 	EMIOENET0TXRRD = 0;
  assign 	EMIOENET0TXRSTATUS = 0;
  assign 	EMIOENET1DMABUSWIDTH = 0;
  assign 	EMIOENET1DMATXENDTOG = 0;
  assign 	EMIOENET1GMIITXD = 0;
  assign 	EMIOENET1GMIITXEN = 0;
  assign 	EMIOENET1GMIITXER = 0;
  assign 	EMIOENET1MDIOMDC = 0;
  assign 	EMIOENET1MDIOO = 0;
  assign 	EMIOENET1MDIOTN = 0;
  assign 	EMIOENET1RXWDATA = 0;
  assign 	EMIOENET1RXWEOP = 0;
  assign 	EMIOENET1RXWERR = 0;
  assign 	EMIOENET1RXWFLUSH = 0;
  assign 	EMIOENET1RXWSOP = 0;
  assign 	EMIOENET1RXWSTATUS = 0;
  assign 	EMIOENET1RXWWR = 0;
  assign 	EMIOENET1SPEEDMODE = 0;
  assign 	EMIOENET1TXRRD = 0;
  assign 	EMIOENET1TXRSTATUS = 0;
  assign 	EMIOGEM0DELAYREQRX = 0;
  assign 	EMIOGEM0DELAYREQTX = 0;
  assign 	EMIOGEM0PDELAYREQRX = 0;
  assign 	EMIOGEM0PDELAYREQTX = 0;
  assign 	EMIOGEM0PDELAYRESPRX = 0;
  assign 	EMIOGEM0PDELAYRESPTX = 0;
  assign 	EMIOGEM0RXSOF = 0;
  assign 	EMIOGEM0SYNCFRAMERX = 0;
  assign 	EMIOGEM0SYNCFRAMETX = 0;
  assign 	EMIOGEM0TSUTIMERCMPVAL = 0;
  assign 	EMIOGEM0TXRFIXEDLAT = 0;
  assign 	EMIOGEM0TXSOF = 0;
  assign 	EMIOGEM1DELAYREQRX = 0;
  assign 	EMIOGEM1DELAYREQTX = 0;
  assign 	EMIOGEM1PDELAYREQRX = 0;
  assign 	EMIOGEM1PDELAYREQTX = 0;
  assign 	EMIOGEM1PDELAYRESPRX = 0;
  assign 	EMIOGEM1PDELAYRESPTX = 0;
  assign 	EMIOGEM1RXSOF = 0;
  assign 	EMIOGEM1SYNCFRAMERX = 0;
  assign 	EMIOGEM1SYNCFRAMETX = 0;
  assign 	EMIOGEM1TSUTIMERCMPVAL = 0;
  assign 	EMIOGEM1TXRFIXEDLAT = 0;
  assign 	EMIOGEM1TXSOF = 0;
  assign   	EMIOGPIO2O = 0;
  assign   	EMIOGPIO2TN = 0;
  assign 	EMIOI2C0SCLO = 0;
  assign 	EMIOI2C0SCLTN = 0;
  assign 	EMIOI2C0SDAO = 0;
  assign 	EMIOI2C0SDATN = 0;
  assign 	EMIOI2C1SCLO = 0;
  assign 	EMIOI2C1SCLTN = 0;
  assign 	EMIOI2C1SDAO = 0;
  assign 	EMIOI2C1SDATN = 0;
  assign 	EMIOSPI0MO = 0;
  assign 	EMIOSPI0MOTN = 0;
  assign 	EMIOSPI0SCLKO = 0;
  assign 	EMIOSPI0SCLKTN = 0;
  assign 	EMIOSPI0SO = 0;
  assign 	EMIOSPI0SSNTN = 0;
  assign   	EMIOSPI0SSON = 0;
  assign 	EMIOSPI0STN = 0;
  assign 	EMIOSPI1MO = 0;
  assign 	EMIOSPI1MOTN = 0;
  assign 	EMIOSPI1SCLKO = 0;
  assign 	EMIOSPI1SCLKTN = 0;
  assign 	EMIOSPI1SO = 0;
  assign 	EMIOSPI1SSNTN = 0;
  assign   	EMIOSPI1SSON = 0;
  assign 	EMIOSPI1STN = 0;
  assign   	EMIOTTC0WAVEO = 0;
  assign   	EMIOTTC1WAVEO = 0;
  assign   	EMIOTTC2WAVEO = 0;
  assign   	EMIOTTC3WAVEO = 0;
  assign 	EMIOU2DSPORTVBUSCTRLUSB30 = 0;
  assign 	FMIOFPDGWDTWS0 = 0;
  assign 	FMIOFPDGWDTWS1 = 0;
  assign   	FMIOFPDLPDEMIOIN = 0;
  assign 	FMIOFPDWWDTINTERRUPT = 0;
  assign 	FMIOFPDWWDTRESET = 0;
  assign 	FMIOFPDWWDTRESETPENDING = 0;
  assign   	FMIOGEM0ADDMATCHVEC = 0;
  assign 	FMIOGEM0RXDATABUFWRQ0 = 0;
  assign 	FMIOGEM0RXDATABUFWRQ1 = 0;
  assign   	FMIOGEM0RXWQUEUE = 0;
  assign   	FMIOGEM0TXRQUEUE = 0;
  assign   	FMIOGEM0TXRTIMESTAMP = 0;
  assign   	FMIOGEM1ADDMATCHVEC = 0;
  assign 	FMIOGEM1RXDATABUFWRQ0 = 0;
  assign 	FMIOGEM1RXDATABUFWRQ1 = 0;
  assign   	FMIOGEM1RXWQUEUE = 0;
  assign   	FMIOGEM1TXRQUEUE = 0;
  assign   	FMIOGEM1TXRTIMESTAMP = 0;
  assign   	FMIOGPIOOEN = 0;
  assign   	FMIOGPIOOUT = 0;
  assign 	FMIOGWDTWS0 = 0;
  assign 	FMIOGWDTWS1 = 0;
  assign 	FMIOI2CSCLOEN = 0;
  assign 	FMIOI2CSCLOUT = 0;
  assign 	FMIOI2CSDAOEN = 0;
  assign 	FMIOI2CSDAOUT = 0;
  assign   	FMIOLPDPMCEMIOIN = 0;
  assign 	FMIOSD0BUSPOWEROUT = 0;
  assign   	FMIOSD0BUSVOLTAGEOUT = 0;
  assign 	FMIOSD0DLLTESTCLK0 = 0;
  assign 	FMIOSD0DLLTESTCLKRX = 0;
  assign 	FMIOSD0DLLTESTCLKTX = 0;
  assign   	FMIOSD0DLLTESTOUT = 0;
  assign 	FMIOSD0LEDCONTROLOUT = 0;
  assign 	FMIOSD0SDIFCLKOUT = 0;
  assign 	FMIOSD0SDIFCMDOE = 0;
  assign 	FMIOSD0SDIFCMDOUT = 0;
  assign   	FMIOSD0SDIFDATOE = 0;
  assign   	FMIOSD0SDIFDATOUT = 0;
  assign 	FMIOSD1BUSPOWEROUT = 0;
  assign   	FMIOSD1BUSVOLTAGEOUT = 0;
  assign 	FMIOSD1DLLTESTCLK0 = 0;
  assign 	FMIOSD1DLLTESTCLKRX = 0;
  assign 	FMIOSD1DLLTESTCLKTX = 0;
  assign   	FMIOSD1DLLTESTOUT = 0;
  assign 	FMIOSD1LEDCONTROLOUT = 0;
  assign 	FMIOSD1SDIFCLKOUT = 0;
  assign 	FMIOSD1SDIFCMDOE = 0;
  assign 	FMIOSD1SDIFCMDOUT = 0;
  assign   	FMIOSD1SDIFDATOE = 0;
  assign   	FMIOSD1SDIFDATOUT = 0;
  assign 	FMIOSYSMONI2CSCLTRIB = 0;
  assign 	FMIOSYSMONI2CSDATRIB = 0;
  assign 	FMIOSYSMONI2CSMBALERTTRIB = 0;
  assign 	FMIOUART0NSIROUT = 0;
  assign 	FMIOUART0NUARTDTR = 0;
  assign 	FMIOUART0NUARTOUT1 = 0;
  assign 	FMIOUART0NUARTOUT2 = 0;
  assign 	FMIOUART0NUARTRTS = 0;
  assign 	FMIOUART0TXD = 0;
  assign 	FMIOUART1NSIROUT = 0;
  assign 	FMIOUART1NUARTDTR = 0;
  assign 	FMIOUART1NUARTOUT1 = 0;
  assign 	FMIOUART1NUARTOUT2 = 0;
  assign 	FMIOUART1NUARTRTS = 0;
  assign 	FMIOUART1TXD = 0;
  assign 	FMIOWWDTINTERRUPT = 0;
  assign 	FMIOWWDTRESET = 0;
  assign 	FMIOWWDTRESETPENDING = 0;
  assign	IFPMCCFUSEUCFUSEUCRCERROR = 0;
  assign 	IFPMCCFUSEUCFUSEUECCERROR = 0;
  assign 	IFPMCCFUSEUCFUSEUENDOFCALIB = 0;
  assign 	IFPMCCFUSEUCFUSEUHALTED = 0;
  assign 	IFPMCCFUSEUCFUSEUHEARTBEAT = 0;
  assign   	IFPSCPMCHANNEL0XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL0XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL0XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL0XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL10XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL10XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL10XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL10XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL11XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL11XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL11XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL11XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL12XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL12XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL12XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL12XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL13XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL13XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL13XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL13XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL14XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL14XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL14XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL14XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL15XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL15XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL15XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL15XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL1XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL1XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL1XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL1XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL2XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL2XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL2XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL2XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL3XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL3XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL3XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL3XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL4XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL4XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL4XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL4XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL5XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL5XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL5XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL5XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL6XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL6XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL6XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL6XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL7XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL7XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL7XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL7XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL8XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL8XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL8XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL8XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMCHANNEL9XPIPEPOWERDOWN = 0;
  assign   	IFPSCPMCHANNEL9XPIPERXPOLARITY = 0;
  assign   	IFPSCPMCHANNEL9XPIPERXTERMINATION = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXCHARISK = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXCOMPLIANCE = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXDATA = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXDATAVALID = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXDEEMPH = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXDETECTRXLOOPBACK = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXELECIDLE = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXMAINCURSOR = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXMARGIN = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXPOSTCURSOR = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXPRECURSOR = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXSTARTBLOCK = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXSWING = 0;
  assign   	IFPSCPMCHANNEL9XPIPETXSYNCHEADER = 0;
  assign   	IFPSCPMHSDPCHANNEL0XPIPERXGEARBOXSLIP = 0;
  assign   	IFPSCPMHSDPCHANNEL0XPIPERXPCSRESET = 0;
  assign   	IFPSCPMHSDPCHANNEL0XPIPETXHEADER = 0;
  assign   	IFPSCPMHSDPCHANNEL0XPIPETXSEQUENCE = 0;
  assign   	IFPSCPMHSDPCHANNEL1XPIPERXGEARBOXSLIP = 0;
  assign   	IFPSCPMHSDPCHANNEL1XPIPERXPCSRESET = 0;
  assign   	IFPSCPMHSDPCHANNEL1XPIPETXHEADER = 0;
  assign   	IFPSCPMHSDPCHANNEL1XPIPETXSEQUENCE = 0;
  assign   	IFPSCPMHSDPCHANNEL2XPIPERXGEARBOXSLIP = 0;
  assign   	IFPSCPMHSDPCHANNEL2XPIPERXPCSRESET = 0;
  assign   	IFPSCPMHSDPCHANNEL2XPIPETXHEADER = 0;
  assign   	IFPSCPMHSDPCHANNEL2XPIPETXSEQUENCE = 0;
  assign   	IFPSCPMHSDPLINKXPIPEGTRXUSRCLK = 0;
  assign   	IFPSCPMINTQUADXPIPEPHYREADYFRBOT = 0;
  assign   	IFPSCPMLINK0XPIPEGTPIPECLK = 0;
  assign   	IFPSCPMLINK0XPIPEPCIELINKREACHTARGET = 0;
  assign   	IFPSCPMLINK0XPIPEPCIELTSSMSTATE = 0;
  assign   	IFPSCPMLINK0XPIPEPCIEPERSTN = 0;
  assign   	IFPSCPMLINK0XPIPEPHYESMADAPTATIONSAVE = 0;
  assign   	IFPSCPMLINK0XPIPEPIPERATE = 0;
  assign   	IFPSCPMLINK1XPIPEGTPIPECLK = 0;
  assign   	IFPSCPMLINK1XPIPEPCIELINKREACHTARGET = 0;
  assign   	IFPSCPMLINK1XPIPEPCIELTSSMSTATE = 0;
  assign   	IFPSCPMLINK1XPIPEPCIEPERSTN = 0;
  assign   	IFPSCPMLINK1XPIPEPHYESMADAPTATIONSAVE = 0;
  assign   	IFPSCPMLINK1XPIPEPIPERATE = 0;
  assign   	IFPSCPMPCSRECOECO = 0;
  assign   	IFPSCPMPCSRPCRAPBEN = 0;
  assign   	IFPSCPMPCSRPCRDISNPICLK = 0;
  assign   	IFPSCPMPCSRPCRFABRICEN = 0;
  assign   	IFPSCPMPCSRPCRGATEREG = 0;
  assign   	IFPSCPMPCSRPCRHOLDSTATE = 0;
  assign   	IFPSCPMPCSRPCRINITSTATE = 0;
  assign   	IFPSCPMPCSRPCRMEMCLR = 0;
  assign   	IFPSCPMPCSRPCRODISABLE = 0;
  assign   	IFPSCPMPCSRPCRPCOMPLETE = 0;
  assign   	IFPSCPMPCSRPCRPWRDN = 0;
  assign   	IFPSCPMPCSRPCRSCANCLR = 0;
  assign   	IFPSCPMPCSRPCRSTARTBISR = 0;
  assign   	IFPSCPMPCSRPCRSTARTCAL = 0;
  assign   	IFPSCPMPCSRPCRTRISTATE = 0;
  assign   	IFPSCPMQUAD0XPIPERXMARGINREQCMD = 0;
  assign   	IFPSCPMQUAD0XPIPERXMARGINREQLANENUM = 0;
  assign   	IFPSCPMQUAD0XPIPERXMARGINREQPAYLOAD = 0;
  assign   	IFPSCPMQUAD0XPIPERXMARGINREQREQ = 0;
  assign   	IFPSCPMQUAD0XPIPERXMARGINRESACK = 0;
  assign   	IFPSCPMQUAD1XPIPERXMARGINREQCMD = 0;
  assign   	IFPSCPMQUAD1XPIPERXMARGINREQLANENUM = 0;
  assign   	IFPSCPMQUAD1XPIPERXMARGINREQPAYLOAD = 0;
  assign   	IFPSCPMQUAD1XPIPERXMARGINREQREQ = 0;
  assign   	IFPSCPMQUAD1XPIPERXMARGINRESACK = 0;
  assign   	IFPSCPMQUAD2XPIPERXMARGINREQCMD = 0;
  assign   	IFPSCPMQUAD2XPIPERXMARGINREQLANENUM = 0;
  assign   	IFPSCPMQUAD2XPIPERXMARGINREQPAYLOAD = 0;
  assign   	IFPSCPMQUAD2XPIPERXMARGINREQREQ = 0;
  assign   	IFPSCPMQUAD2XPIPERXMARGINRESACK = 0;
  assign   	IFPSCPMQUAD3XPIPERXMARGINREQCMD = 0;
  assign   	IFPSCPMQUAD3XPIPERXMARGINREQLANENUM = 0;
  assign   	IFPSCPMQUAD3XPIPERXMARGINREQPAYLOAD = 0;
  assign   	IFPSCPMQUAD3XPIPERXMARGINREQREQ = 0;
  assign   	IFPSCPMQUAD3XPIPERXMARGINRESACK = 0;
  assign   	IFPSOCM2APBPADDR = 0;
  assign   	IFPSOCM2APBPENABLE = 0;
  assign   	IFPSOCM2APBPPROT = 0;
  assign   	IFPSOCM2APBPSEL = 0;
  assign   	IFPSOCM2APBPSTRB = 0;
  assign   	IFPSOCM2APBPWDATA = 0;
  assign   	IFPSOCM2APBPWRITE = 0;
  assign   	IFSYSMONROOTUSERMUXADDR = 0;
  assign   	LPDCPMSWITCHTIMEOUTCNT = 0;
  assign   	LPDRCLKCLK = 0;
  assign   	NCI_NOC_0 = 0;
  assign   	NCI_NOC_1 = 0;
  assign   	NPICLK = 0;
  assign   	NPIRSTN = 0;
  assign   	OSCRTCCLK = 0;
  assign   	PCIE_NOC_0 = 0;
  assign   	PCIE_NOC_1 = 0;
  assign   	PERST0N = 0;
  assign   	PERST1N = 0;
  assign   	PLHSDPEGRESSTDATA = 0;
  assign   	PLHSDPEGRESSTKEEP = 0;
  assign   	PLHSDPEGRESSTLAST = 0;
  assign   	PLHSDPEGRESSTUSER = 0;
  assign   	PLHSDPEGRESSTVALID = 0;
  assign   	PLHSDPINGRESSTREADY = 0;
  assign   	PLPSSMMUARREADY = 0;
  assign   	PLPSSMMUAWREADY = 0;
  assign   	PLPSSMMUCOMPRDREADY = 0;
  assign   	PLPSSMMUCOMPWRREADY = 0;
  assign   	PLREFCLKMUXMONITOR = 0;
  //assign   	PLRST0N = 0;
  //assign   	PLRST1N = 0;
  //assign   	PLRST2N = 0;
  //assign   	PLRST3N = 0;
  assign   	PMCERRORTOPL = 0;
  assign   	PMCPLGPO = 0;
  assign   	PMCPLSYSMONROOTALARM = 0;
  assign   	PMCPLSYSMONROOTNEWDATA = 0;
  //assign   	PMCRCLKCLK = 0;
  assign   	PMC_NOC_0 = 0;
  assign   	PMUAIBAFIFMFPDREQ = 0;
  assign   	PMUAIBAFIFMLPDREQ = 0;
  assign   	PMUERRORTOPL = 0;
  assign   	PSMERRORTOPL = 0;
  assign   	PSPLAFVALID = 0;
  assign   	PSPLATREADY = 0;
  assign   	PSPLEVENTO = 0;
  assign   	PSPLSTANDBYWFE = 0;
  assign   	PSPLSTANDBYWFI = 0;
  assign   	PSPLSYNCREQ = 0;
  assign   	PSPLTRACECTL = 0;
  assign   	PSPLTRACEDATA = 0;
  assign   	PSPLTRIGACK = 0;
  assign   	PSPLTRIGGER = 0;
  assign   	PSSMMUPLARADDR = 0;
  assign   	PSSMMUPLARCACHE = 0;
  assign   	PSSMMUPLARID = 0;
  assign   	PSSMMUPLARVALID = 0;
  assign   	PSSMMUPLAWADDR = 0;
  assign   	PSSMMUPLAWCACHE = 0;
  assign   	PSSMMUPLAWID = 0;
  assign   	PSSMMUPLAWVALID = 0;
  assign   	PSSMMUPLBID = 0;
  assign   	PSSMMUPLBRESP = 0;
  assign   	PSSMMUPLBVALID = 0;
  assign   	PSSMMUPLRERR = 0;
  assign   	PSSMMUPLRID = 0;
  assign   	PSSMMUPLRNS = 0;
  assign   	PSSMMUPLRRESP = 0;
  assign   	PSSMMUPLRVALID = 0;
  assign   	PSSMMUPLWERR = 0;
  assign   	PSSMMUPLWNS = 0;
  assign   	RPUEVENTO0 = 0;
  assign   	RPUEVENTO1 = 0;
  assign   	RPU_NOC_0 = 0;
  assign   	SACEFPDACADDR = 0;
  assign   	SACEFPDACPROT = 0;
  assign   	SACEFPDACSNOOP = 0;
  assign   	SACEFPDACVALID = 0;
  assign   	SACEFPDCDREADY = 0;
  assign   	SACEFPDCRREADY = 0;
  assign   	SAXIGP2RACOUNT = 0;
  assign   	SAXIGP2RCOUNT = 0;
  assign   	SAXIGP2WACOUNT = 0;
  assign   	SAXIGP2WCOUNT = 0;
  assign   	SAXIGP0WACOUNT = 0;
  assign   	SAXIGP0WCOUNT = 0;
  assign   	SAXIGP4RACOUNT = 0;
  assign   	SAXIGP4RCOUNT = 0;
  assign   	SAXIGP4WACOUNT = 0;
  assign   	SAXIGP4WCOUNT = 0;
  assign   	USRCAPTURE = 0;
  assign   	USRDRCK = 0;
  assign   	USRRESET = 0;
  assign   	USRRUNTEST = 0;
  assign   	USRSEL = 0;
  assign   	USRSHIFT = 0;
  assign   	USRTCK = 0;
  assign   	USRTDI = 0;
  assign   	USRTMS = 0;
  assign   	USRUPDATE = 0;


////////////////////////Everest Unused Ports////////////////////////////
//
///* ------------------------------------------- */
///* MIO */
///* ------------------------------------------- */
//
//   always@(PSS_ALTO_CORE_PAD_MIO)
//   begin
//     if(PSS_ALTO_CORE_PAD_MIO !== 0)
//     $display("[%0d] : %0s : MIO is not supported.",$time, DISP_ERR);
//   end
//   
//   assign EMIOCAN0PHYTX = 0;
//   assign EMIOCAN1PHYTX = 0;
//   always @(EMIOCAN0PHYRX or EMIOCAN1PHYRX)
//   begin 
//    if(EMIOCAN0PHYRX | EMIOCAN1PHYRX)
//     $display("[%0d] : %0s : CAN Interface is not supported.",$time, DISP_ERR);
//   end
//
//
//   always @(EMIOENETTSUCLK or
//            EMIOENET0GMIICOL or
//            EMIOENET0GMIICRS or
//            EMIOENET0GMIIRXCLK or
//            EMIOENET0GMIIRXD or
//            EMIOENET0GMIIRXDV or
//            EMIOENET0GMIIRXER or
//            EMIOENET0GMIITXCLK or
//            EMIOENET0MDIOI or
//            EMIOENET0RXWOVERFLOW or
//            EMIOENET0TXRCONTROL or
//            EMIOENET0TXRDATA or
//            EMIOENET0TXRDATARDY or
//            EMIOENET0TXREOP or
//            EMIOENET0TXRERR or
//            EMIOENET0TXRFLUSHED or
//            EMIOENET0TXRSOP or
//            EMIOENET0TXRUNDERFLOW or
//            EMIOENET0TXRVALID or
//            EMIOGEM0TSUINCCTRL)
//    begin
//	  if (EMIOENETTSUCLK |
//          EMIOENET0GMIICOL |
//          EMIOENET0GMIICRS |
//          EMIOENET0GMIIRXCLK |
//          EMIOENET0GMIIRXD |
//          EMIOENET0GMIIRXDV |
//          EMIOENET0GMIIRXER |
//          EMIOENET0GMIITXCLK |
//          EMIOENET0MDIOI |
//          EMIOENET0RXWOVERFLOW |
//          EMIOENET0TXRCONTROL |
//          EMIOENET0TXRDATA |
//          EMIOENET0TXRDATARDY |
//          EMIOENET0TXREOP |
//          EMIOENET0TXRERR |
//          EMIOENET0TXRFLUSHED |
//          EMIOENET0TXRSOP |
//          EMIOENET0TXRUNDERFLOW |
//          EMIOENET0TXRVALID |
//          EMIOGEM0TSUINCCTRL)
//        $display("[%0d] : %0s : GEM Interface is not supported.",$time, DISP_ERR);
//	end
//
//   assign EMIOENET0DMABUSWIDTH = 0;
//   assign EMIOENET0DMATXENDTOG = 0;
//   assign EMIOENET0GEMTSUTIMERCNT = 0;
//   assign EMIOENET0GMIITXD = 0;
//   assign EMIOENET0GMIITXEN = 0;
//   assign EMIOENET0GMIITXER = 0;
//   assign EMIOENET0MDIOMDC = 0;
//   assign EMIOENET0MDIOO = 0;
//   assign EMIOENET0MDIOTN = 0;
//   assign EMIOENET0RXWDATA = 0;
//   assign EMIOENET0RXWEOP = 0;
//   assign EMIOENET0RXWERR = 0;
//   assign EMIOENET0RXWFLUSH = 0;
//   assign EMIOENET0RXWSOP = 0;
//   assign EMIOENET0RXWSTATUS = 0;
//   assign EMIOENET0RXWWR = 0;
//   assign EMIOENET0SPEEDMODE = 0;
//   assign EMIOENET0TXRRD = 0;
//   assign EMIOENET0TXRSTATUS = 0;
//   assign EMIOGEM0DELAYREQRX = 0;
//   assign EMIOGEM0DELAYREQTX = 0;
//   assign EMIOGEM0PDELAYREQRX = 0;
//   assign EMIOGEM0PDELAYREQTX = 0;
//   assign EMIOGEM0PDELAYRESPRX = 0;
//   assign EMIOGEM0PDELAYRESPTX = 0;
//   assign EMIOGEM0RXSOF = 0;
//   assign EMIOGEM0SYNCFRAMERX = 0;
//   assign EMIOGEM0SYNCFRAMETX = 0;
//   assign EMIOGEM0TSUTIMERCMPVAL = 0;
//   assign EMIOGEM0TXRFIXEDLAT = 0;
//   assign EMIOGEM0TXSOF = 0;
//
//   always @(EMIOENETTSUCLK or
//            EMIOENET1GMIICOL or
//            EMIOENET1GMIICRS or
//            EMIOENET1GMIIRXCLK or
//            EMIOENET1GMIIRXD or
//            EMIOENET1GMIIRXDV or
//            EMIOENET1GMIIRXER or
//            EMIOENET1GMIITXCLK or
//            EMIOENET1MDIOI or
//            EMIOENET1RXWOVERFLOW or
//            EMIOENET1TXRCONTROL or
//            EMIOENET1TXRDATA or
//            EMIOENET1TXRDATARDY or
//            EMIOENET1TXREOP or
//            EMIOENET1TXRERR or
//            EMIOENET1TXRFLUSHED or
//            EMIOENET1TXRSOP or
//            EMIOENET1TXRUNDERFLOW or
//            EMIOENET1TXRVALID or
//            EMIOGEM1TSUINCCTRL)
//    begin
//	  if (EMIOENETTSUCLK |
//          EMIOENET1GMIICOL |
//          EMIOENET1GMIICRS |
//          EMIOENET1GMIIRXCLK |
//          EMIOENET1GMIIRXD |
//          EMIOENET1GMIIRXDV |
//          EMIOENET1GMIIRXER |
//          EMIOENET1GMIITXCLK |
//          EMIOENET1MDIOI |
//          EMIOENET1RXWOVERFLOW |
//          EMIOENET1TXRCONTROL |
//          EMIOENET1TXRDATA |
//          EMIOENET1TXRDATARDY |
//          EMIOENET1TXREOP |
//          EMIOENET1TXRERR |
//          EMIOENET1TXRFLUSHED |
//          EMIOENET1TXRSOP |
//          EMIOENET1TXRUNDERFLOW |
//          EMIOENET1TXRVALID |
//          EMIOGEM1TSUINCCTRL)
//        $display("[%0d] : %0s : GEM Interface is not supported.",$time, DISP_ERR);
//	end
//
//   assign EMIOENET1DMABUSWIDTH = 0;
//   assign EMIOENET1DMATXENDTOG = 0;
//   assign EMIOENET1GMIITXD = 0;
//   assign EMIOENET1GMIITXEN = 0;
//   assign EMIOENET1GMIITXER = 0;
//   assign EMIOENET1MDIOMDC = 0;
//   assign EMIOENET1MDIOMDCINT = 0;
//   assign EMIOENET1MDIOO = 0;
//   assign EMIOENET1MDIOTN = 0;
//   assign EMIOENET1RXWDATA = 0;
//   assign EMIOENET1RXWEOP = 0;
//   assign EMIOENET1RXWERR = 0;
//   assign EMIOENET1RXWFLUSH = 0;
//   assign EMIOENET1RXWSOP = 0;
//   assign EMIOENET1RXWSTATUS = 0;
//   assign EMIOENET1RXWWR = 0;
//   assign EMIOENET1SPEEDMODE = 0;
//   assign EMIOENET1TXRRD = 0;
//   assign EMIOENET1TXRSTATUS = 0;
//   assign EMIOGEM1DELAYREQRX = 0;
//   assign EMIOGEM1DELAYREQTX = 0;
//   assign EMIOGEM1PDELAYREQRX = 0;
//   assign EMIOGEM1PDELAYREQTX = 0;
//   assign EMIOGEM1PDELAYRESPRX = 0;
//   assign EMIOGEM1PDELAYRESPTX = 0;
//   assign EMIOGEM1RXSOF = 0;
//   assign EMIOGEM1SYNCFRAMERX = 0;
//   assign EMIOGEM1SYNCFRAMETX = 0;
//   assign EMIOGEM1TSUTIMERCMPVAL = 0;
//   assign EMIOGEM1TXRFIXEDLAT = 0;
//   assign EMIOGEM1TXSOF = 0;
//   assign EMIOGPIO2O = 0;
//   assign EMIOGPIO2TN = 0;
//
//   always @(EMIOENETTSUCLK or
//            EMIOENET2GMIICOL or
//            EMIOENET2GMIICRS or
//            EMIOENET2GMIIRXCLK or
//            EMIOENET2GMIIRXD or
//            EMIOENET2GMIIRXDV or
//            EMIOENET2GMIIRXER or
//            EMIOENET2GMIITXCLK or
//            EMIOENET2MDIOI or
//            EMIOENET2RXWOVERFLOW or
//            EMIOENET2TXRCONTROL or
//            EMIOENET2TXRDATA or
//            EMIOENET2TXRDATARDY or
//            EMIOENET2TXREOP or
//            EMIOENET2TXRERR or
//            EMIOENET2TXRFLUSHED or
//            EMIOENET2TXRSOP or
//            EMIOENET2TXRUNDERFLOW or
//            EMIOENET2TXRVALID or
//            EMIOGEM2TSUINCCTRL)
//    begin
//	  if (EMIOENETTSUCLK |
//          EMIOENET2GMIICOL |
//          EMIOENET2GMIICRS |
//          EMIOENET2GMIIRXCLK |
//          EMIOENET2GMIIRXD |
//          EMIOENET2GMIIRXDV |
//          EMIOENET2GMIIRXER |
//          EMIOENET2GMIITXCLK |
//          EMIOENET2MDIOI |
//          EMIOENET2RXWOVERFLOW |
//          EMIOENET2TXRCONTROL |
//          EMIOENET2TXRDATA |
//          EMIOENET2TXRDATARDY |
//          EMIOENET2TXREOP |
//          EMIOENET2TXRERR |
//          EMIOENET2TXRFLUSHED |
//          EMIOENET2TXRSOP |
//          EMIOENET2TXRUNDERFLOW |
//          EMIOENET2TXRVALID |
//          EMIOGEM2TSUINCCTRL)
//        $display("[%0d] : %0s : GEM Interface is not supported.",$time, DISP_ERR);
//	end
//
//   assign EMIOENET2DMABUSWIDTH = 0;
//   assign EMIOENET2DMATXENDTOG = 0;
//   assign EMIOENET2GMIITXD = 0;
//   assign EMIOENET2GMIITXEN = 0;
//   assign EMIOENET2GMIITXER = 0;
//   assign EMIOENET2MDIOMDC = 0;
//   assign EMIOENET2MDIOO = 0;
//   assign EMIOENET2MDIOTN = 0;
//   assign EMIOENET2RXWDATA = 0;
//   assign EMIOENET2RXWEOP = 0;
//   assign EMIOENET2RXWERR = 0;
//   assign EMIOENET2RXWFLUSH = 0;
//   assign EMIOENET2RXWSOP = 0;
//   assign EMIOENET2RXWSTATUS = 0;
//   assign EMIOENET2RXWWR = 0;
//   assign EMIOENET2SPEEDMODE = 0;
//   assign EMIOENET2TXRRD = 0;
//   assign EMIOENET2TXRSTATUS = 0;
//   assign EMIOGEM2DELAYREQRX = 0;
//   assign EMIOGEM2DELAYREQTX = 0;
//   assign EMIOGEM2PDELAYREQRX = 0;
//   assign EMIOGEM2PDELAYREQTX = 0;
//   assign EMIOGEM2PDELAYRESPRX = 0;
//   assign EMIOGEM2PDELAYRESPTX = 0;
//   assign EMIOGEM2RXSOF = 0;
//   assign EMIOGEM2SYNCFRAMERX = 0;
//   assign EMIOGEM2SYNCFRAMETX = 0;
//   assign EMIOGEM2TSUTIMERCMPVAL = 0;
//   assign EMIOGEM2TXRFIXEDLAT = 0;
//   assign EMIOGEM2TXSOF = 0;
//
//   always @(EMIOENETTSUCLK or
//            EMIOENET3GMIICOL or
//            EMIOENET3GMIICRS or
//            EMIOENET3GMIIRXCLK or
//            EMIOENET3GMIIRXD or
//            EMIOENET3GMIIRXDV or
//            EMIOENET3GMIIRXER or
//            EMIOENET3GMIITXCLK or
//            EMIOENET3MDIOI or
//            EMIOENET3RXWOVERFLOW or
//            EMIOENET3TXRCONTROL or
//            EMIOENET3TXRDATA or
//            EMIOENET3TXRDATARDY or
//            EMIOENET3TXREOP or
//            EMIOENET3TXRERR or
//            EMIOENET3TXRFLUSHED or
//            EMIOENET3TXRSOP or
//            EMIOENET3TXRUNDERFLOW or
//            EMIOENET3TXRVALID or
//            EMIOGEM3TSUINCCTRL)
//    begin
//	  if (EMIOENETTSUCLK |
//          EMIOENET3GMIICOL |
//          EMIOENET3GMIICRS |
//          EMIOENET3GMIIRXCLK |
//          EMIOENET3GMIIRXD |
//          EMIOENET3GMIIRXDV |
//          EMIOENET3GMIIRXER |
//          EMIOENET3GMIITXCLK |
//          EMIOENET3MDIOI |
//          EMIOENET3RXWOVERFLOW |
//          EMIOENET3TXRCONTROL |
//          EMIOENET3TXRDATA |
//          EMIOENET3TXRDATARDY |
//          EMIOENET3TXREOP |
//          EMIOENET3TXRERR |
//          EMIOENET3TXRFLUSHED |
//          EMIOENET3TXRSOP |
//          EMIOENET3TXRUNDERFLOW |
//          EMIOENET3TXRVALID |
//          EMIOGEM3TSUINCCTRL)
//        $display("[%0d] : %0s : GEM Interface is not supported.",$time, DISP_ERR);
//	end
//
//   assign EMIOENET3DMABUSWIDTH = 0;
//   assign EMIOENET3DMATXENDTOG = 0;
//   assign EMIOENET3GMIITXD = 0;
//   assign EMIOENET3GMIITXEN = 0;
//   assign EMIOENET3GMIITXER = 0;
//   assign EMIOENET3MDIOMDC = 0;
//   assign EMIOENET3MDIOO = 0;
//   assign EMIOENET3MDIOTN = 0;
//   assign EMIOENET3RXWDATA = 0;
//   assign EMIOENET3RXWEOP = 0;
//   assign EMIOENET3RXWERR = 0;
//   assign EMIOENET3RXWFLUSH = 0;
//   assign EMIOENET3RXWSOP = 0;
//   assign EMIOENET3RXWSTATUS = 0;
//   assign EMIOENET3RXWWR = 0;
//   assign EMIOENET3SPEEDMODE = 0;
//   assign EMIOENET3TXRRD = 0;
//   assign EMIOENET3TXRSTATUS = 0;
//   assign EMIOGEM3DELAYREQRX = 0;
//   assign EMIOGEM3DELAYREQTX = 0;
//   assign EMIOGEM3PDELAYREQRX = 0;
//   assign EMIOGEM3PDELAYREQTX = 0;
//   assign EMIOGEM3PDELAYRESPRX = 0;
//   assign EMIOGEM3PDELAYRESPTX = 0;
//   assign EMIOGEM3RXSOF = 0;
//   assign EMIOGEM3SYNCFRAMERX = 0;
//   assign EMIOGEM3SYNCFRAMETX = 0;
//   assign EMIOGEM3TSUTIMERCMPVAL = 0;
//   assign EMIOGEM3TXRFIXEDLAT = 0;
//   assign EMIOGEM3TXSOF = 0;
//
//   always @(EMIOGPIOI)
//     begin
//	   if(EMIOGPIOI)
//        $display("[%0d] : %0s : GPIO Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOGPIOO = 0;
//   assign EMIOGPIOTN = 0;
//
//   always @(EMIOHUBPORTOVERCRNTUSB20 or
//            EMIOHUBPORTOVERCRNTUSB21 or
//            EMIOHUBPORTOVERCRNTUSB30 or
//            EMIOHUBPORTOVERCRNTUSB31 or
//            EMIOU2DSPORTVBUSCTRLUSB30 or 
//            EMIOU2DSPORTVBUSCTRLUSB31 or
//            EMIOU3DSPORTVBUSCTRLUSB30 or
//            EMIOU3DSPORTVBUSCTRLUSB31)
//     begin
//	   if(EMIOHUBPORTOVERCRNTUSB20 |
//          EMIOHUBPORTOVERCRNTUSB21 |
//          EMIOHUBPORTOVERCRNTUSB30 |
//          EMIOHUBPORTOVERCRNTUSB31 |
//		  EMIOU2DSPORTVBUSCTRLUSB30 | 
//          EMIOU2DSPORTVBUSCTRLUSB31 |
//          EMIOU3DSPORTVBUSCTRLUSB30 |
//          EMIOU3DSPORTVBUSCTRLUSB31)
//         $display("[%0d] : %0s : USB Interface is not supported.",$time, DISP_ERR);
//	 end
//	
//    always @(EMIOI2C0SCLI or
//             EMIOI2C0SDAI or
//             EMIOI2C1SCLI or
//             EMIOI2C1SDAI)
//	  begin
//        if(EMIOI2C0SCLI |
//           EMIOI2C0SDAI |
//           EMIOI2C1SCLI |
//           EMIOI2C1SDAI)
//         $display("[%0d] : %0s : I2C Interface is not supported.",$time, DISP_ERR);
//	  end
//
//   assign EMIOI2C0SCLO = 0;
//   assign EMIOI2C0SCLTN = 0;
//   assign EMIOI2C0SDAO = 0;
//   assign EMIOI2C0SDATN = 0;
//   assign EMIOI2C1SCLO = 0;
//   assign EMIOI2C1SCLTN = 0;
//   assign EMIOI2C1SDAO = 0;
//   assign EMIOI2C1SDATN = 0;
//
//   always @(EMIOSDIO0CDN or
//            EMIOSDIO0CMDIN or
//            EMIOSDIO0DATAIN or
//            EMIOSDIO0FBCLKIN or
//            EMIOSDIO0WP or
//            EMIOSDIO1CDN or
//            EMIOSDIO1CMDIN or
//            EMIOSDIO1DATAIN or
//            EMIOSDIO1FBCLKIN or
//            EMIOSDIO1WP)
//     begin
//	   if(EMIOSDIO0CDN |
//          EMIOSDIO0CMDIN |
//          EMIOSDIO0DATAIN |
//          EMIOSDIO0FBCLKIN |
//          EMIOSDIO0WP |
//          EMIOSDIO1CDN |
//          EMIOSDIO1CMDIN |
//          EMIOSDIO1DATAIN |
//          EMIOSDIO1FBCLKIN |
//          EMIOSDIO1WP)
//         $display("[%0d] : %0s : SDIO Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOSDIO0BUSPOWER = 0;
//   assign EMIOSDIO0BUSVOLT = 0;
//   assign EMIOSDIO0CLKOUT = 0;
//   assign EMIOSDIO0CMDENA = 0;
//   assign EMIOSDIO0CMDOUT = 0;
//   assign EMIOSDIO0DATAENA = 0;
//   assign EMIOSDIO0DATAOUT = 0;
//   assign EMIOSDIO0LEDCONTROL = 0;
//   assign EMIOSDIO1BUSPOWER = 0;
//   assign EMIOSDIO1BUSVOLT = 0;
//   assign EMIOSDIO1CLKOUT = 0;
//   assign EMIOSDIO1CMDENA = 0;
//   assign EMIOSDIO1CMDOUT = 0;
//   assign EMIOSDIO1DATAENA = 0;
//   assign EMIOSDIO1DATAOUT = 0;
//   assign EMIOSDIO1LEDCONTROL = 0;
//
//   always @(EMIOSPI0MI or
//            EMIOSPI0SCLKI or
//            EMIOSPI0SI or
//            EMIOSPI0SSIN or
//            EMIOSPI1MI or
//            EMIOSPI1SCLKI or
//            EMIOSPI1SI or
//            EMIOSPI1SSIN)
//     begin
//      if(EMIOSPI0MI |
//         EMIOSPI0SCLKI |
//         EMIOSPI0SI |
//         EMIOSPI0SSIN |
//         EMIOSPI1MI |
//         EMIOSPI1SCLKI |
//         EMIOSPI1SI |
//         EMIOSPI1SSIN)
//        $display("[%0d] : %0s : SPI Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOSPI0MO = 0;
//   assign EMIOSPI0MOTN = 0;
//   assign EMIOSPI0SCLKO = 0;
//   assign EMIOSPI0SCLKOINT = 0;
//   assign EMIOSPI0SCLKTN = 0;
//   assign EMIOSPI0SO = 0;
//   assign EMIOSPI0SSNTN = 0;
//   assign EMIOSPI0SSON = 0;
//   assign EMIOSPI0STN = 0;
//   assign EMIOSPI1MO = 0;
//   assign EMIOSPI1MOTN = 0;
//   assign EMIOSPI1SCLKO = 0;
//   assign EMIOSPI1SCLKTN = 0;
//   assign EMIOSPI1SO = 0;
//   assign EMIOSPI1SSNTN = 0;
//   assign EMIOSPI1SSON = 0;
//   assign EMIOSPI1STN = 0;
//
//   always @(EMIOTTC0CLKI or
//            EMIOTTC1CLKI or
//            EMIOTTC2CLKI or
//            EMIOTTC3CLKI)
//     begin
//	   if(EMIOTTC0CLKI |
//          EMIOTTC1CLKI |
//          EMIOTTC2CLKI |
//          EMIOTTC3CLKI)
//        $display("[%0d] : %0s : TTC Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOTTC0WAVEO = 0;
//   assign EMIOTTC1WAVEO = 0;
//   assign EMIOTTC2WAVEO = 0;
//   assign EMIOTTC3WAVEO = 0;
//
//   always @(EMIOUART0CTSN or
//            EMIOUART0DCDN or
//            EMIOUART0DSRN or
//            EMIOUART0RIN or
//            EMIOUART0RX or
//            EMIOUART1CTSN or
//            EMIOUART1DCDN or
//            EMIOUART1DSRN or
//            EMIOUART1RIN or
//            EMIOUART1RX)
//     begin
//	   if(EMIOUART0CTSN |
//          EMIOUART0DCDN |
//          EMIOUART0DSRN |
//          EMIOUART0RIN |
//          EMIOUART0RX |
//          EMIOUART1CTSN |
//          EMIOUART1DCDN |
//          EMIOUART1DSRN |
//          EMIOUART1RIN |
//          EMIOUART1RX)
//        $display("[%0d] : %0s : TTC Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOUART0DTRN = 0;
//   assign EMIOUART0RTSN = 0;
//   assign EMIOUART0TX = 0;
//   assign EMIOUART1DTRN = 0;
//   assign EMIOUART1RTSN = 0;
//   assign EMIOUART1TX = 0;
//
//   always @(EMIOWDT0CLKI or
//            EMIOWDT1CLKI)
//     begin
//	   if(EMIOWDT0CLKI |
//          EMIOWDT1CLKI)
//        $display("[%0d] : %0s : WDT Interface is not supported.",$time, DISP_ERR);
//	 end
//
//   assign EMIOWDT0RSTO = 0;
//   assign EMIOWDT1RSTO = 0;
//
//   assign ADMA2PLCACK = 0;
//   assign ADMA2PLTVLD = 0;
//   assign CFUEOS = 0;
//   assign CPMOSCCLKDIV2 = 0;
//   assign APLLTESTCLKOUT = 0;
//   assign BSCANTDO = 0;
//   assign DBGPATHFIFOBYPASS = 0;
//   assign DDRDTO = 0;
//   assign DPAUDIOREFCLK = 0;
//   assign DPAUXDATAOEN = 0;
//   assign DPAUXDATAOUT = 0;
//   assign DPLIVEVIDEODEOUT = 0;
//   assign DPLLTESTCLKOUT = 0;
//   assign DPMAXISMIXEDAUDIOTDATA = 0;
//   assign DPMAXISMIXEDAUDIOTID = 0;
//   assign DPMAXISMIXEDAUDIOTVALID = 0;
//   assign DPSAXISAUDIOTREADY = 0;
//   assign DPVIDEOOUTHSYNC = 0;
//   assign DPVIDEOOUTPIXEL1 = 0;
//   assign DPVIDEOOUTVSYNC = 0;
//   assign DPVIDEOREFCLK = 0;
//   assign FMIOFPDGWDTWS0 = 0;
//   assign FMIOFPDGWDTWS1 = 0;
//   assign FMIOFPDLPDEMIOIN = 0;
//   assign FMIOFPDWWDTINTERRUPT = 0;
//   assign FMIOFPDWWDTRESET = 0;
//   assign FMIOFPDWWDTRESETPENDING = 0;
//   assign FMIOGEM0ADDMATCHVEC = 0;
//   assign FMIOGEM0RXDATABUFWRQ0 = 0;
//   assign FMIOGEM0RXDATABUFWRQ1 = 0;
//   assign FMIOGEM0RXWQUEUE = 0;
//   assign FMIOGEM0TXRQUEUE = 0;
//   assign FMIOGEM0TXRTIMESTAMP = 0;
//   assign FMIOGEM1ADDMATCHVEC = 0;
//   assign FMIOGEM1RXDATABUFWRQ0 = 0;
//   assign FMIOGEM1RXDATABUFWRQ1 = 0;
//   assign FMIOGEM1RXWQUEUE = 0;
//   assign FMIOGEM1TXRQUEUE = 0;
//   assign FMIOGEM1TXRTIMESTAMP = 0;
//   assign FMIOGPIOOEN = 0;
//   assign FMIOGPIOOUT = 0;
//   assign FMIOGWDTWS0 = 0;
//   assign FMIOGWDTWS1 = 0;
//   assign FMIOI2CSCLOEN = 0;
//   assign FMIOI2CSCLOUT = 0;
//   assign FMIOI2CSDAOEN = 0;
//   assign FMIOI2CSDAOUT = 0;
//   assign FMIOLPDPMCEMIOIN = 0;
//   assign FMIOSD0BUSPOWEROUT = 0;
//   assign FMIOSD0BUSVOLTAGEOUT = 0;
//   assign FMIOSD0DLLTESTCLK0 = 0;
//   assign FMIOSD0DLLTESTCLKRX = 0;
//   assign FMIOSD0DLLTESTCLKTX = 0;
//   assign FMIOCHARAFIFSFPDTESTOUTPUT = 0;
//   assign FMIOCHARAFIFSLPDTESTOUTPUT = 0;
//   assign FMIOCHARGEMTESTOUTPUT = 0;
//   assign FMIOGEMTSUCLKTOPLBUFG = 0;
//   assign FMIOGEM0FIFORXCLKTOPLBUFG = 0;
//   assign FMIOGEM0FIFOTXCLKTOPLBUFG = 0;
//   assign FMIOGEM1FIFORXCLKTOPLBUFG = 0;
//   assign FMIOGEM1FIFOTXCLKTOPLBUFG = 0;
//   assign FMIOGEM2FIFORXCLKTOPLBUFG = 0;
//   assign FMIOGEM2FIFOTXCLKTOPLBUFG = 0;
//   assign FMIOGEM3FIFORXCLKTOPLBUFG = 0;
//   assign FMIOGEM3FIFOTXCLKTOPLBUFG = 0;
//   assign FMIOSD0DLLTESTOUT = 0;
//   assign FMIOSD0SDIFCMDOUT = 0;
//   assign FMIOSD0SDIFDATOE = 0;
//   assign FMIOSD0SDIFDATOUT = 0;
//   assign FMIOSD1BUSPOWEROUT = 0;
//   assign FMIOSD1BUSVOLTAGEOUT = 0;
//   assign FMIOSD0LEDCONTROLOUT = 0;
//   assign FMIOSD0SDIFCLKOUT = 0;
//   assign FMIOSD1SDIFCLKOUTINT = 0;
//   assign FMIOSD0SDIFCLKOUTINT = 0;
//   assign FMIOSD1SDIFCMDOE = 0;
//   assign FMIOSD0SDIFCMDOE = 0;
//   assign FMIOSD1DLLTESTOUT = 0;
//   assign FMIOSD1SDIFCMDOUT = 0;
//   assign FMIOSD1SDIFDATOE = 0;
//   assign FMIOSD1SDIFDATOUT = 0;
//   assign FMIOSYSMONI2CSCLTRIB = 0;
//   assign FMIOSYSMONI2CSDATRIB = 0;
//   assign FMIOSD1LEDCONTROLOUT = 0;
//   assign FMIOSYSMONI2CSDATRIB = 0;
//   assign FMIOUART0NSIROUT = 0;
//   assign FMIOUART0NUARTDTR = 0;
//   assign FMIOUART0NUARTOUT1 = 0;
//   assign FMIOUART0NUARTOUT2 = 0;
//   assign FMIOUART0NUARTRTS = 0;
//   assign FMIOUART0TXD = 0;
//   assign FMIOUART1TXD = 0;
//   assign FMIOWWDTINTERRUPT = 0;
//   assign FMIOWWDTRESET = 0;
//   assign FMIOWWDTRESETPENDING = 0;
//   assign FMIOUART1NSIROUT = 0;
//   assign FMIOUART1NUARTDTR = 0;
//   assign FMIOUART1NUARTOUT1 = 0;
//   assign FMIOUART1NUARTOUT2 = 0;
//   assign FMIOUART1NUARTRTS = 0;
//   assign FMIOSD1DLLTESTCLK0 = 0;
//   assign FMIOSD1DLLTESTCLKRX = 0;
//   assign FMIOSD1DLLTESTCLKTX = 0;
//   assign FMIOTESTIOCHARSCANOUT = 0;
//   assign FPDPLLTESTOUT = 0;
//   assign FPDPLSPARE0OUT = 0;
//   assign FPDPLSPARE1OUT = 0;
//   assign FPDPLSPARE2OUT = 0;
//   assign FPDPLSPARE3OUT = 0;
//   assign FPDPLSPARE4OUT = 0;
//   assign FTMGPO = 0;
//   assign GDMA2PLCACK = 0;
//   assign GDMA2PLTVLD = 0;
//   assign IOCHARAUDIOOUTTESTDATA = 0;
//   assign IOCHARVIDEOOUTTESTDATA = 0;
//   assign IOPLLTESTCLKOUT = 0;
//
//  assign IFPSCPMCHANNEL0XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL0XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL0XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL0XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL0XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL0XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL0XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL0XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL0XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL10XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL10XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL10XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL10XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL10XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL10XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL10XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL10XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL10XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL11XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL11XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL11XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL11XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL11XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL11XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL11XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL11XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL11XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL12XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL12XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL12XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL12XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL12XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL12XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL12XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL12XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL12XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL13XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL13XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL13XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL13XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL13XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL13XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL13XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL13XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL13XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL14XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL14XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL14XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL14XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL14XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL14XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL14XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL14XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL14XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL15XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL15XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL15XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL15XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL15XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL15XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL15XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL15XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL15XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL1XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL1XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL1XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL1XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL1XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL1XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL1XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL1XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL1XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL2XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL2XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL2XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL2XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL2XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL2XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL2XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL2XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL2XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL3XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL3XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL3XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL3XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL3XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL3XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL3XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL3XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL3XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL4XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL4XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL4XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL4XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL4XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL4XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL4XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL4XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL4XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL5XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL5XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL5XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL5XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL5XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL5XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL5XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL5XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL5XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL6XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL6XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL6XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL6XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL6XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL6XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL6XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL6XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL6XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL7XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL7XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL7XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL7XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL7XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL7XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL7XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL7XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL7XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL8XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL8XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL8XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL8XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL8XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL8XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL8XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL8XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL8XPIPERXVALID = 0;
//  assign IFPSCPMCHANNEL9XPIPEPHYSTATUS = 0;
//  assign IFPSCPMCHANNEL9XPIPERXCHARISK = 0;
//  assign IFPSCPMCHANNEL9XPIPERXDATA = 0;
//  assign IFPSCPMCHANNEL9XPIPERXDATAVALID = 0;
//  assign IFPSCPMCHANNEL9XPIPERXELECIDLE = 0;
//  assign IFPSCPMCHANNEL9XPIPERXSTARTBLOCK = 0;
//  assign IFPSCPMCHANNEL9XPIPERXSTATUS = 0;
//  assign IFPSCPMCHANNEL9XPIPERXSYNCHEADER = 0;
//  assign IFPSCPMCHANNEL9XPIPERXVALID = 0;
//  assign IFPSCPMHSDPCHANNEL0XPIPERXDATAVALID = 0;
//  assign IFPSCPMHSDPCHANNEL0XPIPERXHEADER = 0;
//  assign IFPSCPMHSDPCHANNEL0XPIPERXHEADERVALID = 0;
//  assign IFPSCPMHSDPCHANNEL0XPIPERXRESETDONE = 0;
//  assign IFPSCPMHSDPCHANNEL0XPIPETXRESETDONE = 0;
//  assign IFPSCPMHSDPCHANNEL1XPIPERXDATAVALID = 0;
//  assign IFPSCPMHSDPCHANNEL1XPIPERXHEADER = 0;
//  assign IFPSCPMHSDPCHANNEL1XPIPERXHEADERVALID = 0;
//  assign IFPSCPMHSDPCHANNEL1XPIPERXRESETDONE,
//  IFPSCPMHSDPCHANNEL1XPIPETXRESETDONE = 0;
//  assign IFPSCPMHSDPCHANNEL2XPIPERXDATAVALID = 0;
//  assign IFPSCPMHSDPCHANNEL2XPIPERXHEADER = 0;
//  assign IFPSCPMHSDPCHANNEL2XPIPERXHEADERVALID = 0;
//  assign IFPSCPMHSDPCHANNEL2XPIPERXRESETDONE = 0;
//  assign IFPSCPMHSDPCHANNEL2XPIPETXRESETDONE = 0;
//  assign IFPSCPMHSDPLINKXPIPEGTRXOUTCLK = 0;
//  assign IFPSCPMINTQUADXPIPEPHYREADYTOBOT = 0;
//  assign IFPSCPMLINK0XPIPEBUFGTCE = 0;
//  assign IFPSCPMLINK0XPIPEBUFGTCEMASK = 0;
//  assign IFPSCPMLINK0XPIPEBUFGTDIV = 0;
//  assign IFPSCPMLINK0XPIPEBUFGTRST = 0;
//  assign IFPSCPMLINK0XPIPEBUFGTRSTMASK = 0;
//  assign IFPSCPMLINK0XPIPEGTOUTCLK = 0;
//  assign IFPSCPMLINK0XPIPEPHYREADY = 0;
//  assign IFPSCPMLINK1XPIPEBUFGTCE = 0;
//  assign IFPSCPMLINK1XPIPEBUFGTCEMASK = 0;
//  assign IFPSCPMLINK1XPIPEBUFGTDIV = 0;
//  assign IFPSCPMLINK1XPIPEBUFGTRST = 0;
//  assign IFPSCPMLINK1XPIPEBUFGTRSTMASK = 0;
//  assign IFPSCPMLINK1XPIPEGTOUTCLK = 0;
//  assign IFPSCPMLINK1XPIPEPHYREADY = 0;
//
//  assign IFPSOCM2APBPRDATA = 0;
//  assign IFPSOCM2APBPREADY = 0;
//  assign IFPSOCM2APBPSLVERR = 0;
//
//  assign MJTAGTCK = 0;
//  assign MJTAGTDI = 0;
//  assign MJTAGTMS = 0;
//  assign NFIQ0LPDRPU = 0;
//  assign NFIQ1LPDRPU = 0;
//  assign NIRQ0LPDRPU = 0;
//  assign NIRQ1LPDRPU = 0;
//  assign NPIINTERRUPTOUT = 0;
//  assign PL2ADMACVLD = 0;
//  assign PL2ADMATACK = 0;
//  assign PLACECLK = 0;
//  assign PLACPINACT = 0;
//  assign PLCONFIGDONE = 0;
//  assign PLFPDAUXREFCLK = 0;
//  assign PLHSDPCLK = 0;
//  assign PLHSDPEGRESSTREADY = 0;
//  assign PLHSDPINGRESSTDATA = 0;
//  assign PLHSDPINGRESSTKEEP = 0;
//  assign PLHSDPINGRESSTLAST = 0;
//  assign PLHSDPINGRESSTVALID = 0;
//  assign PLLPDAUXREFCLK = 0;
//  assign PLPMCAUXREFCLK = 0;
//  assign PLPMCFPGACLOCKSTOP = 0;
//  assign PLPSAFREADY = 0;
//  assign PLPSAPUGICFIQ = 0;
//  assign PLPSAPUGICIRQ = 0;
//  assign PLPSATBCLK = 0;
//  assign PLPSATBYTES = 0;
//  assign PLPSATDATA = 0;
//  assign PLPSATID = 0;
//  assign PLPSATVALID = 0;
//  assign PLPSEVENTI = 0;
//  assign PLPSIRQ0 = 0;
//  assign PLPSIRQ1 = 0;
//  assign PLPSSMMUARADDR = 0;
//  assign PLPSSMMUARCACHE = 0;
//  assign PLPSSMMUARID = 0;
//  assign PLPSSMMUARVALID = 0;
//  assign PLPSSMMUAWADDR = 0;
//  assign PLPSSMMUAWCACHE = 0;
//  assign PLPSSMMUAWID = 0;
//  assign PLPSSMMUAWVALID = 0;
//  assign PLPSSMMUCLOCK = 0;
//  assign PLPSSMMUCOMPRDID = 0;
//  assign PLPSSMMUCOMPRDVAL = 0;
//  assign PLPSSMMUCOMPWRID = 0;
//  assign PLPSSMMUCOMPWRVAL = 0;
//  assign PLPSSMMURNS = 0;
//  assign PLPSSMMURSMID = 0;
//  assign PLPSSMMUWNS = 0;
//  assign PLPSSMMUWSMID = 0;
//  assign PLPSTRACECLK = 0;
//  assign PLPSTRIGACK = 0;
//  assign PLPSTRIGGER = 0;
//  assign PMCPLGPI = 0;
//  assign PMCPLIRQ = 0;
//  assign PMUERRORFROMPL = 0;
//  assign PSSMMUPLARREADY = 0;
//  assign PSSMMUPLAWREADY = 0;
//  assign PSSMMUPLBREADY = 0;
//  assign PSSMMUPLRREADY = 0;
//  assign PSS_PAD_RTCPADI = 0;
//  assign RPUEVENTI0 = 0;
//  assign RPUEVENTI1 = 0;
//  assign RTCPADI = 0;
//  assign STMEVENT = 0;
//  assign USRTDO = 0;
//  assign DBGSE = 0;
//
//
//  assign IFPSCPMPCSRPSRBISRDONE = 0;
//  assign IFPSCPMPCSRPSRBISRERR = 0;
//  assign IFPSCPMPCSRPSRCALDONE = 0;
//  assign IFPSCPMPCSRPSRCALERROR = 0;
//  assign IFPSCPMPCSRPSRINCAL = 0;
//  assign IFPSCPMPCSRPSRMEMCLRDONE = 0;
//  assign IFPSCPMPCSRPSRMEMCLRPASS = 0;
//  assign IFPSCPMPCSRPSRSCANCLRDONE = 0;
//  assign IFPSCPMPCSRPSRSCANCLRPASS = 0;
//  assign IFPSCPMQUAD0XPIPERXMARGINREQACK = 0;
//  assign IFPSCPMQUAD0XPIPERXMARGINRESCMD = 0;
//  assign IFPSCPMQUAD0XPIPERXMARGINRESLANENUM = 0;
//  assign IFPSCPMQUAD0XPIPERXMARGINRESPAYLOAD = 0;
//  assign IFPSCPMQUAD0XPIPERXMARGINRESREQ = 0;
//  assign IFPSCPMQUAD1XPIPERXMARGINREQACK = 0;
//  assign IFPSCPMQUAD1XPIPERXMARGINRESCMD = 0;
//  assign IFPSCPMQUAD1XPIPERXMARGINRESLANENUM = 0;
//  assign IFPSCPMQUAD1XPIPERXMARGINRESPAYLOAD = 0;
//  assign IFPSCPMQUAD1XPIPERXMARGINRESREQ = 0;
//  assign IFPSCPMQUAD2XPIPERXMARGINREQACK = 0;
//  assign IFPSCPMQUAD2XPIPERXMARGINRESCMD = 0;
//  assign IFPSCPMQUAD2XPIPERXMARGINRESLANENUM = 0;
//  assign IFPSCPMQUAD2XPIPERXMARGINRESPAYLOAD = 0;
//  assign IFPSCPMQUAD2XPIPERXMARGINRESREQ = 0;
//  assign IFPSCPMQUAD3XPIPERXMARGINREQACK = 0;
//  assign IFPSCPMQUAD3XPIPERXMARGINRESCMD = 0;
//  assign IFPSCPMQUAD3XPIPERXMARGINRESLANENUM = 0;
//  assign IFPSCPMQUAD3XPIPERXMARGINRESPAYLOAD = 0;
//  assign IFPSCPMQUAD3XPIPERXMARGINRESREQ = 0;
//
//
//   assign LPDPLLTESTOUT = 0;
//   assign LPDPLSPARE0OUT = 0;
//   assign LPDPLSPARE1OUT = 0;
//   assign LPDPLSPARE2OUT = 0;
//   assign LPDPLSPARE3OUT = 0;
//   assign LPDPLSPARE4OUT = 0;
//   assign OAFECMNCALIBCOMPOUT = 0;
//   assign OAFEPGAVDDCR = 0;
//   assign OAFEPGAVDDIO = 0;
//   assign OAFEPGDVDDCR = 0;
//   assign OAFEPGSTATICAVDDCR = 0;
//   assign OAFEPGSTATICAVDDIO = 0;
//   assign OAFEPLLCLKSYMHS = 0;
//   assign OAFEPLLDCOCOUNT = 0;
//   assign OAFEPLLFBCLKFRAC = 0;
//   assign OAFERXHSRXCLOCKSTOPACK = 0;
//   assign OAFERXPIPELFPSBCNRXELECIDLE = 0;
//   assign OAFERXPIPESIGDET = 0;
//   assign OAFERXSYMBOL = 0;
//   assign OAFERXSYMBOLCLKBY2 = 0;
//   assign OAFERXUPHYRXCALIBDONE = 0;
//   assign OAFERXUPHYSAVECALCODE = 0;
//   assign OAFERXUPHYSAVECALCODEDATA = 0;
//   assign OAFERXUPHYSTARTLOOPBUF = 0;
//   assign OAFETXDIGRESETRELACK = 0;
//   assign OAFETXPIPETXDNRXDET = 0;
//   assign OAFETXPIPETXDPRXDET = 0;
//   assign ODBGL0PHYSTATUS = 0;
//   assign ODBGL0POWERDOWN = 0;
//   assign ODBGL0RATE = 0;
//   assign ODBGL0RSTB = 0;
//   assign ODBGL0RXCLK = 0;
//   assign ODBGL0RXDATA = 0;
//   assign ODBGL0RXDATAK = 0;
//   assign ODBGL0RXELECIDLE = 0;
//   assign ODBGL0RXPOLARITY = 0;
//   assign ODBGL0RXSGMIIENCDET = 0;
//   assign ODBGL0RXSTATUS = 0;
//   assign ODBGL0RXVALID = 0;
//   assign ODBGL0SATACORECLOCKREADY = 0;
//   assign ODBGL0SATACOREREADY = 0;
//   assign ODBGL0SATACORERXDATA = 0;
//   assign ODBGL0SATACORERXDATAVALID = 0;
//   assign ODBGL0SATACORERXSIGNALDET = 0;
//   assign ODBGL0SATAPHYCTRLPARTIAL = 0;
//   assign ODBGL0SATAPHYCTRLRESET = 0;
//   assign ODBGL0SATAPHYCTRLRXRATE = 0;
//   assign ODBGL0SATAPHYCTRLRXRST = 0;
//   assign ODBGL0SATAPHYCTRLSLUMBER = 0;
//   assign ODBGL0SATAPHYCTRLTXDATA = 0;
//   assign ODBGL0SATAPHYCTRLTXIDLE = 0;
//   assign ODBGL0SATAPHYCTRLTXRATE = 0;
//   assign ODBGL0SATAPHYCTRLTXRST = 0;
//   assign ODBGL0TXCLK = 0;
//   assign ODBGL0TXDATA = 0;
//   assign ODBGL0TXDATAK = 0;
//   assign ODBGL0TXDETRXLPBACK = 0;
//   assign ODBGL0TXELECIDLE = 0;
//   assign ODBGL0TXSGMIIEWRAP = 0;
//   assign ODBGL1PHYSTATUS = 0;
//   assign ODBGL1POWERDOWN = 0;
//   assign ODBGL1RATE = 0;
//   assign ODBGL1RSTB = 0;
//   assign ODBGL1RXCLK = 0;
//   assign ODBGL1RXDATA = 0;
//   assign ODBGL1RXDATAK = 0;
//   assign ODBGL1RXELECIDLE = 0;
//   assign ODBGL1RXPOLARITY = 0;
//   assign ODBGL1RXSGMIIENCDET = 0;
//   assign ODBGL1RXSTATUS = 0;
//   assign ODBGL1RXVALID = 0;
//   assign ODBGL1SATACORECLOCKREADY = 0;
//   assign ODBGL1SATACOREREADY = 0;
//   assign ODBGL1SATACORERXDATA = 0;
//   assign ODBGL1SATACORERXDATAVALID = 0;
//   assign ODBGL1SATACORERXSIGNALDET = 0;
//   assign ODBGL1SATAPHYCTRLPARTIAL = 0;
//   assign ODBGL1SATAPHYCTRLRESET = 0;
//   assign ODBGL1SATAPHYCTRLRXRATE = 0;
//   assign ODBGL1SATAPHYCTRLRXRST = 0;
//   assign ODBGL1SATAPHYCTRLSLUMBER = 0;
//   assign ODBGL1SATAPHYCTRLTXDATA = 0;
//   assign ODBGL1SATAPHYCTRLTXIDLE = 0;
//   assign ODBGL1SATAPHYCTRLTXRATE = 0;
//   assign ODBGL1SATAPHYCTRLTXRST = 0;
//   assign ODBGL1TXCLK = 0;
//   assign ODBGL1TXDATA = 0;
//   assign ODBGL1TXDATAK = 0;
//   assign ODBGL1TXDETRXLPBACK = 0;
//   assign ODBGL1TXELECIDLE = 0;
//   assign ODBGL1TXSGMIIEWRAP = 0;
//   assign ODBGL2PHYSTATUS = 0;
//   assign ODBGL2POWERDOWN = 0;
//   assign ODBGL2RATE = 0;
//   assign ODBGL2RSTB = 0;
//   assign ODBGL2RXCLK = 0;
//   assign ODBGL2RXDATA = 0;
//   assign ODBGL2RXDATAK = 0;
//   assign ODBGL2RXELECIDLE = 0;
//   assign ODBGL2RXPOLARITY = 0;
//   assign ODBGL2RXSGMIIENCDET = 0;
//   assign ODBGL2RXSTATUS = 0;
//   assign ODBGL2RXVALID = 0;
//   assign ODBGL2SATACORECLOCKREADY = 0;
//   assign ODBGL2SATACOREREADY = 0;
//   assign ODBGL2SATACORERXDATA = 0;
//   assign ODBGL2SATACORERXDATAVALID = 0;
//   assign ODBGL2SATACORERXSIGNALDET = 0;
//   assign ODBGL2SATAPHYCTRLPARTIAL = 0;
//   assign ODBGL2SATAPHYCTRLRESET = 0;
//   assign ODBGL2SATAPHYCTRLRXRATE = 0;
//   assign ODBGL2SATAPHYCTRLRXRST = 0;
//   assign ODBGL2SATAPHYCTRLSLUMBER = 0;
//   assign ODBGL2SATAPHYCTRLTXDATA = 0;
//   assign ODBGL2SATAPHYCTRLTXIDLE = 0;
//   assign ODBGL2SATAPHYCTRLTXRATE = 0;
//   assign ODBGL2SATAPHYCTRLTXRST = 0;
//   assign ODBGL2TXCLK = 0;
//   assign ODBGL2TXDATA = 0;
//   assign ODBGL2TXDATAK = 0;
//   assign ODBGL2TXDETRXLPBACK = 0;
//   assign ODBGL2TXELECIDLE = 0;
//   assign ODBGL2TXSGMIIEWRAP = 0;
//   assign ODBGL3PHYSTATUS = 0;
//   assign ODBGL3POWERDOWN = 0;
//   assign ODBGL3RATE = 0;
//   assign ODBGL3RSTB = 0;
//   assign ODBGL3RXCLK = 0;
//   assign ODBGL3RXDATA = 0;
//   assign ODBGL3RXDATAK = 0;
//   assign ODBGL3RXELECIDLE = 0;
//   assign ODBGL3RXPOLARITY = 0;
//   assign ODBGL3RXSGMIIENCDET = 0;
//   assign ODBGL3RXSTATUS = 0;
//   assign ODBGL3RXVALID = 0;
//   assign ODBGL3SATACORECLOCKREADY = 0;
//   assign ODBGL3SATACOREREADY = 0;
//   assign ODBGL3SATACORERXDATA = 0;
//   assign ODBGL3SATACORERXDATAVALID = 0;
//   assign ODBGL3SATACORERXSIGNALDET = 0;
//   assign ODBGL3SATAPHYCTRLPARTIAL = 0;
//   assign ODBGL3SATAPHYCTRLRESET = 0;
//   assign ODBGL3SATAPHYCTRLRXRATE = 0;
//   assign ODBGL3SATAPHYCTRLRXRST = 0;
//   assign ODBGL3SATAPHYCTRLSLUMBER = 0;
//   assign ODBGL3SATAPHYCTRLTXDATA = 0;
//   assign ODBGL3SATAPHYCTRLTXIDLE = 0;
//   assign ODBGL3SATAPHYCTRLTXRATE = 0;
//   assign ODBGL3SATAPHYCTRLTXRST = 0;
//   assign ODBGL3TXCLK = 0;
//   assign ODBGL3TXDATA = 0;
//   assign ODBGL3TXDATAK = 0;
//   assign ODBGL3TXDETRXLPBACK = 0;
//   assign ODBGL3TXELECIDLE = 0;
//   assign ODBGL3TXSGMIIEWRAP = 0;
//   assign OSCRTCCLK = 0;
//   assign PCAPCSB = 0;
//   assign PCAPPR = 0;
//   assign PCAPRDWRB = 0;
//   assign PCAPWDATA = 0;
//   assign PCAPWDATACLK = 0;
//   assign PCFGBOOT = 0;
//   assign PCFGGSR = 0;
//   assign PCFGGTS = 0;
//   assign PCFGINITB = 0;
//   assign PCFGJTAGCFGDISABLE = 0;
//   assign PCFGPORCNT4K = 0;
//   assign PCFGPROG = 0;
//   assign PCFGTCK = 0;
//   assign PCFGTDI = 0;
//   assign PCFGTMS = 0;
//   assign PMUAIBAFIFMFPDREQ = 0;
//   assign PMUAIBAFIFMLPDREQ = 0;
//   assign PMUERRORTOPL = 0;
//   assign PMUPLGPO = 0;
//   assign PSDADDR = 0;
//   assign PSDCLK = 0;
//   assign PSDEN = 0;
//   assign PSDI = 0;
//   assign PSDWE = 0;
//   assign PSPLEVENTO = 0;
//   assign PSPLIRQFPD = 0;
//   assign PSPLIRQLPD = 0;
//   assign PSPLSTANDBYWFE = 0;
//   assign PSPLSTANDBYWFI = 0;
//   assign PSPLSYSOSCCLK = 0;
//   assign PSPLTRACECTL = 0;
//   assign PSPLTRACEDATA = 0;
//   assign PSPLTRIGACK = 0;
//   assign PSPLTRIGGER = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXN0OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXN1OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXN2OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXN3OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXP0OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXP1OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXP2OUT = 0;
//   assign PSS_ALTO_CORE_PAD_MGTTXP3OUT = 0;
//   assign PSS_ALTO_CORE_PAD_PADO = 0;
//   assign PSTPPLOUT = 0;
//   assign RPLLTESTCLKOUT = 0;
//   assign RPUEVENTO0 = 0;
//   assign RPUEVENTO1 = 0;
//   assign SACEFPDACADDR = 0;
//   assign SACEFPDACPROT = 0;
//   assign SACEFPDACSNOOP = 0;
//   assign SACEFPDACVALID = 0;
//   assign SACEFPDCDREADY = 0;
//   assign SACEFPDCRREADY = 0;
//   assign SYSMONSENSEFULLVCCPSAUXN = 0;
//   assign SYSMONSENSEFULLVCCPSAUXP = 0;
//   assign SYSMONSENSEFULLVCCPSINTFPN = 0;
//   assign SYSMONSENSEFULLVCCPSINTFPP = 0;
//   assign SYSMONSENSEFULLVCCPSINTLPN = 0;
//   assign SYSMONSENSEFULLVCCPSINTLPP = 0;
//   assign TESTADCOUT = 0;
//   assign TESTAMSOSC = 0;
//   assign TESTBSCANTDO = 0;
//   assign TESTDB = 0;
//   assign TESTDDR2PLDCDSKEWOUT = 0;
//   assign TESTDO = 0;
//   assign TESTDRDY = 0;
//   assign TESTMONDATA = 0;
//   assign TESTPLPLLLOCKOUT = 0;
//   assign TESTPLSCANCHOPPERSO = 0;
//   assign TESTPLSCANEDTOUTAPU = 0;
//   assign TESTPLSCANEDTOUTCPU0 = 0;
//   assign TESTPLSCANEDTOUTCPU1 = 0;
//   assign TESTPLSCANEDTOUTCPU2 = 0;
//   assign TESTPLSCANEDTOUTCPU3 = 0;
//   assign TESTPLSCANEDTOUTDDR = 0;
//   assign TESTPLSCANEDTOUTFP = 0;
//   assign TESTPLSCANEDTOUTGPU = 0;
//   assign TESTPLSCANEDTOUTLP = 0;
//   assign TESTPLSCANEDTOUTUSB3 = 0;
//   assign TESTPLSCANSLCRCONFIGSO = 0;
//   assign TESTPLSCANSPAREOUT0 = 0;
//   assign TESTPLSCANSPAREOUT1 = 0;
//   assign TSTRTCCALIBREGOUT = 0;
//   assign TSTRTCOSCCLKOUT = 0;
//   assign TSTRTCOSCCNTRLOUT = 0;
//   assign TSTRTCSECCOUNTEROUT = 0;
//   assign TSTRTCSECONDSRAWINT = 0;
//   assign TSTRTCTICKCOUNTEROUT = 0;
//   assign TSTRTCTIMESETREGOUT = 0;
//   assign UNUSEDTIEHIGH = 0;
//   assign UNUSEDTIELOW = 0;
//   assign VCUPCFGFUSEVCUDISBOT = 0;
//   assign VCUPCFGFUSEVCUDISTOP = 0;
//   assign VPLLTESTCLKOU = 0;
