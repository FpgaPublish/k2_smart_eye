interface data_interface;

logic    [31:0] data;
    
endinterface //data_interface